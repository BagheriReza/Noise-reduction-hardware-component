
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.all;
	USE IEEE.STD_LOGIC_UNSIGNED.all;
ENTITY mux_2to1_nbit IS
	GENERIC(CONSTANT n : INTEGER := 17);
	PORT(sel : IN STD_LOGIC;a,b : IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);c : OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0));
END mux_2to1_nbit;

ARCHITECTURE dataflow OF mux_2to1_nbit IS
BEGIN
c <= a WHEN sel ='1' ELSE b;
END dataflow;